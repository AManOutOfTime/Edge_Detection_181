library verilog;
use verilog.vl_types.all;
entity blur_tb is
end blur_tb;
