library verilog;
use verilog.vl_types.all;
entity sobel_conv_tb is
end sobel_conv_tb;
