library verilog;
use verilog.vl_types.all;
entity sobel_conv_tb2 is
end sobel_conv_tb2;
