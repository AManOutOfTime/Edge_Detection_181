library verilog;
use verilog.vl_types.all;
entity sqrt_approx_tb is
end sqrt_approx_tb;
